// `include "ctrl_encode_def.v"

//123
module ctrl (
    Op,
    Funct7,
    Funct3,
    Zero,
    RegWrite,
    MemWrite,
    EXTOp,
    ALUOp,
    NPCOp,
    ALUSrc,
    GPRSel,
    WDSel,
    DMType
);

  input [6:0] Op;  // opcode
  input [6:0] Funct7;  // funct7
  input [2:0] Funct3;  // funct3
  input Zero;

  output RegWrite;  // control signal for register write
  output MemWrite;  // control signal for memory write
  output [5:0] EXTOp;  // control signal to signed extension
  output [4:0] ALUOp;  // ALU opertion
  output [2:0] NPCOp;  // next pc operation
  output ALUSrc;  // ALU source for A
  output [2:0] DMType;
  output [1:0] GPRSel;  // general purpose register selection
  output [1:0] WDSel;  // (register) write data selection

  // r format
  wire rtype = ~Op[6] & Op[5] & Op[4] & ~Op[3] & ~Op[2] & Op[1] & Op[0];  //0110011
  wire i_add  = rtype& ~Funct7[6]&~Funct7[5]&~Funct7[4]&~Funct7[3]&~Funct7[2]&~Funct7[1]&~Funct7[0]&~Funct3[2]&~Funct3[1]&~Funct3[0]; // add 0000000 000
  wire i_sub  = rtype& ~Funct7[6]& Funct7[5]&~Funct7[4]&~Funct7[3]&~Funct7[2]&~Funct7[1]&~Funct7[0]&~Funct3[2]&~Funct3[1]&~Funct3[0]; // sub 0100000 000
  wire i_or   = rtype& ~Funct7[6]&~Funct7[5]&~Funct7[4]&~Funct7[3]&~Funct7[2]&~Funct7[1]&~Funct7[0]& Funct3[2]& Funct3[1]&~Funct3[0]; // or 0000000 110
  wire i_and  = rtype& ~Funct7[6]&~Funct7[5]&~Funct7[4]&~Funct7[3]&~Funct7[2]&~Funct7[1]&~Funct7[0]& Funct3[2]& Funct3[1]& Funct3[0]; // and 0000000 111


  // i format
  wire itype_l = ~Op[6] & ~Op[5] & ~Op[4] & ~Op[3] & ~Op[2] & Op[1] & Op[0];  //0000011

  wire lw = itype_l & (Funct3 == 3'b010);
  wire lb = itype_l & (Funct3 == 3'b000);
  wire lh = itype_l & (Funct3 == 3'b001);
  wire lbu = itype_l & (Funct3 == 3'b100);
  wire lhu = itype_l & (Funct3 == 3'b101);

  // i format
  wire itype_r = ~Op[6] & ~Op[5] & Op[4] & ~Op[3] & ~Op[2] & Op[1] & Op[0];  //0010011
  wire i_addi = itype_r & ~Funct3[2] & ~Funct3[1] & ~Funct3[0];  // addi 000
  wire i_ori = itype_r & Funct3[2] & Funct3[1] & ~Funct3[0];  // ori 110
  wire i_andi = itype_r & (Funct3 == 3'b111);
  wire i_xori = itype_r & (Funct3 == 3'b100);
  wire i_srai = itype_r & (Funct3 == 3'b101);
  wire i_slli = itype_r & (Funct3 == 3'b001);

  wire lui = (Op == 7'b0110111);
  wire auipc = (Op == 7'b0010111);
  //jalr
  wire i_jalr = Op[6] & Op[5] & ~Op[4] & ~Op[3] & Op[2] & Op[1] & Op[0];  //jalr 1100111

  // s format
  wire stype = ~Op[6] & Op[5] & ~Op[4] & ~Op[3] & ~Op[2] & Op[1] & Op[0];  //0100011
  wire i_sw = stype & ~Funct3[2] & Funct3[1] & ~Funct3[0];  // sw 010

  wire sw = stype & (Funct3 == 3'b010);
  wire sb = stype & (Funct3 == 3'b000);
  wire sh = stype & (Funct3 == 3'b001);

  // sb format
  wire sbtype = Op[6] & Op[5] & ~Op[4] & ~Op[3] & ~Op[2] & Op[1] & Op[0];  //1100011
  wire i_beq = sbtype & ~Funct3[2] & ~Funct3[1] & ~Funct3[0];  // beq

  // j format
  wire i_jal = Op[6] & Op[5] & ~Op[4] & Op[3] & Op[2] & Op[1] & Op[0];  // jal 1101111

  // generate control signals
  assign RegWrite = rtype | itype_r | i_jalr | i_jal | lui | auipc;  // register write
  assign MemWrite = stype;  // memory write
  assign ALUSrc   = itype_r | stype | i_jal | i_jalr | lui | auipc;  // ALU B is from instruction immediate

  // signed extension
  // EXT_CTRL_ITYPE_SHAMT 6'b100000
  // EXT_CTRL_ITYPE	      6'b010000
  // EXT_CTRL_STYPE	      6'b001000
  // EXT_CTRL_BTYPE	      6'b000100
  // EXT_CTRL_UTYPE	      6'b000010
  // EXT_CTRL_JTYPE	      6'b000001
  assign EXTOp[5] = 0;
  //assign EXTOp[4]    =  i_ori | i_andi | i_jalr;
  assign EXTOp[4] = i_ori | i_addi;
  assign EXTOp[3] = stype;
  assign EXTOp[2] = sbtype;
  assign EXTOp[1] = lui | auipc;
  assign EXTOp[0] = i_jal;




  // WDSel_FromALU 2'b00
  // WDSel_FromMEM 2'b01
  // WDSel_FromPC  2'b10 
  assign WDSel[0] = itype_l;
  assign WDSel[1] = i_jal | i_jalr;

  // NPC_PLUS4   3'b000
  // NPC_BRANCH  3'b001
  // NPC_JUMP    3'b010
  // NPC_JALR	3'b100
  assign NPCOp[0] = sbtype & Zero;
  assign NPCOp[1] = i_jal;
  assign NPCOp[2] = i_jalr;



  assign ALUOp[0] = itype_l | stype | i_addi | i_ori | i_add | i_or | lui;
  assign ALUOp[1] = i_jalr | itype_l | stype | i_addi | i_add | i_and | auipc;
  assign ALUOp[2] = i_andi|i_and|i_ori|i_or|i_beq|i_sub;
  assign ALUOp[3] = i_andi|i_and|i_ori|i_or;
  assign ALUOp[4] = 0;

  assign DMType[0] = lh | sh | sb | lb;
  assign DMType[1] = lhu | sb | lb;
  assign DMType[2] = lbu;

endmodule
